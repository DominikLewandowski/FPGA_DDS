`ifndef CONFIG_VH
`define CONFIG_VH

// ------ ROM ------ //
`define ROM_PHASE_MAX_VAL   14'd10000       // Ilo�� pr�bek sygna�u
`define ROM_PHASE_BIT       14              // Ilo�� bit�w potrzebna na zapis fazy

`endif
