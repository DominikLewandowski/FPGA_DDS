`ifndef CONFIG_VH
`define CONFIG_VH

`endif